`timescale 1ns / 1ps

module ro1(
				input en,
				output out
			);
	 
       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5, w6, w7, w8, w9,w10,w11,w12,w13,w14,w15,w16,w17, 
		w18, w19,w20,w21,w22,w23,w24,w25,w26,w27,w28,w29,w30,
		 w31,w32,w33,w34,w35,w36,w37,w38,w39,w40,w41,
       w42, w43,w44,w45, w46, w47, w48, w49,w50 ,
		  w51, w52, w53,w54,w55, w56, w57, w58, w59,w60,
		 w61, w62, w63,w64,w65, w66, w67, w68, w69,w70,
		 w71, w72, w73,w74,w75, w76, w77, w78, w79,w80,
		  w81, w82, w83,w84,w85, w86, w87, w88, w89,w90,
		  w91, w92, w93,w94,w95, w96, w97, w98, w99,w100,
		 w101, w102, w103,w104,w105, w106, w107, w108, w109,w110,
		  w111, w112, w113,w114,w115, w116, w117, w118, w119,w120,
		  w121, w122, w123,w124,w125, w126, w127, w128, w129,w130,
		  w131, w132, w133,w134,w135, w136, w137, w138, w139,w140, w141;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #5(w5, w4);
        not #1(w6, w5);
        not #1(w7, w6);
        not #1(w8, w7);
        not #1(w9, w8);
        not #1(w10, w9);
        not #1(w11, w10);
        not #1(w12, w11);
        not #1(w13, w12);
		  
       not #1(w14, w13);
        not #1(w15, w14);
        not #1(w16, w15);
        not #1(w17, w16);
        not #1(w18, w17);
        not #1(w19, w18);
        not #1(w20, w19);
        not #1(w21, w20);
        not #1(w22, w21);
        not #1(w23, w22);
        not #1(w24, w23);
        not #1(w25, w24);
        not #1(w26, w25);
        not #1(w27, w26);
        not #1(w28, w27);
        not #1(w29, w28);
        not #1(w30, w29);
        not #1(w31, w30);
        not #1(w32, w31);
        not #1(w33, w32);
        not #1(w34, w33);
        not #1(w35, w34);
        not #1(w36, w35);
        not #1(w37, w36);
        not #1(w38, w37);
        not #1(w39, w38);
        not #1(w40, w39);
        not #1(w41, w40);
		  not #1(w42, w41);
		 
        not #1(w43, w42);
        not #1(w44,w43);
        not #1(w45, w44);
        not #1(w46, w45);
        not #1(w47, w46);
        not #1(w48, w47);
        not #1(w49, w48);
        not #1(w50, w49);
		  not #1(w51, w50);
		  not #1(w52, w51);
        not #1(w53, w52);
        not #1(w54, w53);
        not #1(w55, w54);
        not #1(w56, w55);
        not #1(w57, w56);
        not #1(w58, w57);
        not #1(w59, w58);
        not #1(w60, w59);
		  not #1(w61, w60);
		  not #1(w62, w61);
        not #1(w63, w62);
        not #1(w64, w63);
        not #1(w65, w64);
        not #1(w66, w65);
        not #1(w67, w66);
        not #1(w68, w67);
        not #1(w69, w68);
        not #1(w70, w69);
        not #1(w71, w70);
		  
		  not #1(w72, w71);
        not #1(w73, w72);
        not #1(w74, w73);
        not #1(w75, w74);
        not #1(w76, w75);
        not #1(w77, w76);
        not #1(w78, w77);
        not #1(w79, w78);
        not #1(w80, w79);
        not #1(w81, w80);
		  
		  not #1(w82, w81);
        not #1(w83, w82);
        not #1(w84, w83);
        not #1(w85, w84);
        not #1(w86, w85);
        not #1(w87, w86);
        not #1(w88, w87);
        not #1(w89, w88);
        not #1(w90, w89);
        not #1(w91, w90);
		  
		  not #1(w92, w91);
        not #1(w93, w92);
        not #1(w94, w93);
        not #1(w95, w94);
        not #1(w96, w95);
        not #1(w97, w96);
        not #1(w98, w97);
        not #1(w99, w98);
        not #1(w100, w99);
        not #1(w101, w100);
		  
		  not #1(w102, w101);
        not #1(w103, w102);
        not #1(w104, w103);
        not #1(w105, w104);
        not #1(w106, w105);
        not #1(w107, w106);
        not #1(w108, w107);
        not #1(w109, w108);
        not #1(w110, w109);
        not #1(w111, w110);
		  
		  not #1(w112, w111);
        not #1(w113, w112);
        not #1(w114, w113);
        not #1(w115, w114);
        not #1(w116, w115);
        not #1(w117, w116);
        not #1(w118, w117);
        not #1(w119, w118);
        not #1(w120, w119);
        not #1(w121, w120);
		  
		  not #1(w122, w121);
        not #1(w123, w122);
        not #1(w124, w123);
        not #1(w125, w124);
        not #1(w126, w125);
        not #1(w127, w126);
        not #1(w128, w127);
        not #1(w129, w128);
        not #1(w130, w129);
        not #1(w131, w130);
		  
        not #1(w132, w131);
        not #1(w133, w132);
        not #1(w134, w133);
        not #1(w135, w134);
        not #1(w136, w135);
        not #1(w137, w136);
        not #1(w138, w137);
        not #1(w139, w138);
        not #1(w140, w139);
        not #1(w141, w140);
		  
		   not #1(out, w141);
		
endmodule
