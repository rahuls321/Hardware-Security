`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:11:01 08/07/2017 
// Design Name: 
// Module Name:    mux_4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mux_4(input W0,W1,W2,W3,input[1:0] S,output [15:0] M);
wire [15:0] W0,W1,W2,W3;
	
	 assign M[0] = W0[0] & ~S[1] & ~S[0] | W1[0] & ~S[1] & S[0] | W2[0] & S[1] & ~S[0] | W3[0] & S[1] & S[0];
	 assign M[1] = W0[1] & ~S[1] & ~S[0] | W1[1] & ~S[1] & S[0] | W2[1] & S[1] & ~S[0] | W3[1] & S[1] & S[0];
    assign M[2] = W0[2] & ~S[1] & ~S[0] | W1[2] & ~S[1] & S[0] | W2[2] & S[1] & ~S[0] | W3[2] & S[1] & S[0];
    assign M[3] = W0[3] & ~S[1] & ~S[0] | W1[3] & ~S[1] & S[0] | W2[3] & S[1] & ~S[0] | W3[3] & S[1] & S[0];
    assign M[4] = W0[4] & ~S[1] & ~S[0] | W1[4] & ~S[1] & S[0] | W2[4] & S[1] & ~S[0] | W3[4] & S[1] & S[0];
    assign M[5] = W0[5] & ~S[1] & ~S[0] | W1[5] & ~S[1] & S[0] | W2[5] & S[1] & ~S[0] | W3[5] & S[1] & S[0];
    assign M[6] = W0[6] & ~S[1] & ~S[0] | W1[6] & ~S[1] & S[0] | W2[6] & S[1] & ~S[0] | W3[6] & S[1] & S[0];
    assign M[7] = W0[7] & ~S[1] & ~S[0] | W1[7] & ~S[1] & S[0] | W2[7] & S[1] & ~S[0] | W3[7] & S[1] & S[0];
    assign M[8] = W0[8] & ~S[1] & ~S[0] | W1[8] & ~S[1] & S[0] | W2[8] & S[1] & ~S[0] | W3[8] & S[1] & S[0];
	 assign M[9] = W0[9] & ~S[1] & ~S[0] | W1[9] & ~S[1] & S[0] | W2[9] & S[1] & ~S[0] | W3[9] & S[1] & S[0];
    assign M[10] = W0[10] & ~S[1] & ~S[0] | W1[10] & ~S[1] & S[0] | W2[10] & S[1] & ~S[0] | W3[10] & S[1] & S[0];
    assign M[11] = W0[11] & ~S[1] & ~S[0] | W1[11] & ~S[1] & S[0] | W2[11] & S[1] & ~S[0] | W3[11] & S[1] & S[0];
    assign M[12] = W0[12] & ~S[1] & ~S[0] | W1[12] & ~S[1] & S[0] | W2[12] & S[1] & ~S[0] | W3[12] & S[1] & S[0];
    assign M[13] = W0[13] & ~S[1] & ~S[0] | W1[13] & ~S[1] & S[0] | W2[13] & S[1] & ~S[0] | W3[13] & S[1] & S[0];
    assign M[14] = W0[14] & ~S[1] & ~S[0] | W1[14] & ~S[1] & S[0] | W2[14] & S[1] & ~S[0] | W3[14] & S[1] & S[0];
    assign M[15] = W0[15] & ~S[1] & ~S[0] | W1[15] & ~S[1] & S[0] | W2[15] & S[1] & ~S[0] | W3[15] & S[1] & S[0];
	/* assign M[16] = W[16] & ~S[1] & ~S[0] | X[16] & ~S[1] & S[0] | Y[16] & S[1] & ~S[0] | Z[16] & S[1] & S[0];
	 assign M[17] = W[17] & ~S[1] & ~S[0] | X[17] & ~S[1] & S[0] | Y[17] & S[1] & ~S[0] | Z[17] & S[1] & S[0];
    assign M[18] = W[18] & ~S[1] & ~S[0] | X[18] & ~S[1] & S[0] | Y[18] & S[1] & ~S[0] | Z[16] & S[1] & S[0];
    assign M[19] = W[19] & ~S[1] & ~S[0] | X[19] & ~S[1] & S[0] | Y[19] & S[1] & ~S[0] | Z[19] & S[1] & S[0];
    assign M[20] = W[20] & ~S[1] & ~S[0] | X[20] & ~S[1] & S[0] | Y[20] & S[1] & ~S[0] | Z[20] & S[1] & S[0];
    assign M[21] = W[21] & ~S[1] & ~S[0] | X[21] & ~S[1] & S[0] | Y[21] & S[1] & ~S[0] | Z[21] & S[1] & S[0];
    assign M[22] = W[22] & ~S[1] & ~S[0] | X[22] & ~S[1] & S[0] | Y[22] & S[1] & ~S[0] | Z[22] & S[1] & S[0];
    assign M[23] = W[23] & ~S[1] & ~S[0] | X[23] & ~S[1] & S[0] | Y[23] & S[1] & ~S[0] | Z[23] & S[1] & S[0];
    assign M[24] = W[24] & ~S[1] & ~S[0] | X[24] & ~S[1] & S[0] | Y[24] & S[1] & ~S[0] | Z[24] & S[1] & S[0];
	 assign M[25] = W[25] & ~S[1] & ~S[0] | X[25] & ~S[1] & S[0] | Y[25] & S[1] & ~S[0] | Z[25] & S[1] & S[0];
    assign M[26] = W[26] & ~S[1] & ~S[0] | X[26] & ~S[1] & S[0] | Y[26] & S[1] & ~S[0] | Z[26] & S[1] & S[0];
    assign M[27] = W[27] & ~S[1] & ~S[0] | X[27] & ~S[1] & S[0] | Y[27] & S[1] & ~S[0] | Z[27] & S[1] & S[0];
    assign M[28] = W[28] & ~S[1] & ~S[0] | X[28] & ~S[1] & S[0] | Y[28] & S[1] & ~S[0] | Z[28] & S[1] & S[0];
    assign M[29] = W[29] & ~S[1] & ~S[0] | X[29] & ~S[1] & S[0] | Y[29] & S[1] & ~S[0] | Z[29] & S[1] & S[0];
    assign M[30] = W[30] & ~S[1] & ~S[0] | X[30] & ~S[1] & S[0] | Y[30] & S[1] & ~S[0] | Z[30] & S[1] & S[0];
    assign M[31] = W[31] & ~S[1] & ~S[0] | X[31] & ~S[1] & S[0] | Y[31] & S[1] & ~S[0] | Z[31] & S[1] & S[0];
	 
*/
	 endmodule
